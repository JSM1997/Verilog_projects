`include "p_f_module_c_inicial_i_d.v"
`include "p_f_module_c_tipica_i_d.v"
`include "p_f_module_c_final_i_d.v"

module red_izq_der (

    input wire [2:0] palabraA,
    input wire [2:0] palabraB,
    output wire resultado
);



)

endmodule
