module Celda_inicial_d_i #(
    parameter N=3/*preguntar al profe si esta es una definición valida porque no se puede pedir */ 
    
) (/*Celda inicial no tiene entradas de estado presente(son evaluadas), tiene entradas primarias, y salidas de proximo estado*/
    input wire a_p, 
    input wire b_p,
    output wire p_x,
    output wire p_y
);
assing p_x = 
    
endmodule